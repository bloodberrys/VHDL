--LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--USE NUMERIC_STD.ALL;
--
--ENTITY INPUTAN IS
--PORT ( ADDRESSSIGNAL : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
--		 CLOCK : IN STD_LOGIC;
--		 WRITEENABLER : IN STD_LOGIC;
--		 DATA
--		 );
--END COUNTER;
--
--ARCHITECTURE COUNTING OF COUNTER IS
--SIGNAL PENGHITUNG : INTEGER RANGE 0 TO 99;
--BEGIN
--	LOOPING : 
--	for I in 0 RANGE TO 5 loop
--			ADDRESSSIGNAL <= STD_LOGIC_VECTOR(UNSIGNED(ADDRESSSIGNAL + 1));
--	end loop;
--
--END ARCHITECTURE;