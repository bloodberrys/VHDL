LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY SEG7 IS
PORT ( ENABLER : IN STD_LOGIC;
		 NILAI : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 KELUAR : OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END ENTITY;

ARCHITECTURE SEV OF SEG7 IS
BEGIN
PROCESS (NILAI)
BEGIN
CASE NILAI IS
		WHEN "0000" => KELUAR <= "0000000";
		WHEN "0001" => KELUAR <= "0110000";
		WHEN "0010" => KELUAR <= "1101101";
		WHEN "0011" => KELUAR <= "1111001";
		WHEN "0100" => KELUAR <= "0110011";
		WHEN "0101" => KELUAR <= "1011011";
		WHEN "0110" => KELUAR <= "1011111";
		WHEN "0111" => KELUAR <= "1110000";
		WHEN "1000" => KELUAR <= "1111111";
		WHEN "1001" => KELUAR <= "1111011";
		WHEN OTHERS => KELUAR <= "0000000";
END CASE;
END PROCESS;
END ARCHITECTURE;
