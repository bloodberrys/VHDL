LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY COUNTER IS
PORT ( ENABLER : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 CLOCK : IN STD_LOGIC;
		 ANGKA : IN INTEGER RANGE -2 TO 256;
		 OUTPUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COUNTER;

ARCHITECTURE COUNTING OF COUNTER IS
SIGNAL PENGHITUNG : INTEGER RANGE 0 TO 256;
SIGNAL DUMMY : INTEGER RANGE -4 TO 256 := 60;
BEGIN

	PROCESS (clOCK,reset,enabler)
	BEGIN
		if reSET ='1' and enabler ='1' then
					DUMMY <= ANGKA - 1;
					PENGHITUNG <= ANGKA + (((angka /10)*6));
		else
		if RISING_EDGE(CLOCK) THEN
			IF (enabler = '1' and reset ='0' ) THEN
				DUMMY <= DUMMY - 1;
				if DUMMY >= 10 then
				PENGHITUNG <= DUMMY + ((DUMMY / 10)* 6);
				elsif DUMMY < 0 then
				penghitung <= 0;
				else
				penghitung <= DUMMY;
				end if;
			END IF;
		end if;
				OUTPUT <= STD_LOGIC_VECTOR(UNSIGNED(TO_UNSIGNED(PENGHITUNG,8)));
		END IF;
	END PROCESS;
END ARCHITECTURE;