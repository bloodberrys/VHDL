LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DFLIP_FLOP IS
PORT
(

D : IN STD_LOGIC;
CLK : IN STD_LOGIC;
Q,QNOT : OUT STD_LOGIC);
END ENTITY;

ARCHITECTURE DFLIP_FLOP OF DFLIP_FLOP IS
SIGNAL PRESENT : STD_LOGIC;
BEGIN
RISING :PROCESS (CLK,d) IS
BEGIN
if rising_edge(CLK) THEN
	PRESENT <= D;
END IF;
END PROCESS;
Q <= PRESENT;
QNOT <= NOT(PRESENT);
END ARCHITECTURE;
